module debug_var_display_controller(
    input sys_clk,
    input sys_rst_n,
    input [3:0] debug_var,
    input [3:0] debug_var_on,
    output reg [3:0] debug_var_rgb
);





endmodule