module tb_character;




endmodule